PK   WlKTzײ�+*  ��    cirkitFile.json�ێ�F��_��Uy��<��N�
;��a5轐� �RbK�5�Y�nz�ucTVF��g�o�F��I��[~47��O���=6���������t�p�{G�������9��}��pw�~����|�q����<���`�ǡ�ۇ�f?8��PzC�M���T#u�i�n,cƾ�۽ݽ���7�[ ��'1�Ԃ�;1�Ԃ�{1�Ԃ�1�Ԃ��d�}��Ӈ����y_����X�ڏ�	m�Mg���f(��v{W�d�Q�_�}(�`��?<�<<����}.A����y�{���~��_N%v�Ԃ��b���*��ި�I�d���tONx�C� $<H>z�M$
��!6�(d#H)�M�B�1Dl"QHG�#$GH>��M$
�P"6����������%N>��M$
�X�c���%N>��M$
�X"6�(�ɜ�&,�mb
�x�	��&,�b���ꓻ��PX)��{+�|���l@�Ro�G#��D!�%6�( ϲ�#��� b�B>��M$�B���t�'$�R�d@�g|�W�(_9�7���D��k!�	��� b�B>��M$
�"6�(�0_�xNR+%H�0_���f8[�I�!G�&�\��M$
��H�Dl"Q�G�	��V����K��$$�W�#��gk�{C>��M$
��Hr%&6�(�#��D��� b�B>��M$
�"6�(�#�؄�r"6�(�Dl"Q�s�����Ȧ��><<!���&3GK�������.�f�("���c��1(a���a}簾�����=�w�;(a�~��.`}�#,]��`}�����.�1��+��������]���n�-��!K)��TX�WX�C�Kg�5�w5�wP:�����5Xa���߽����&hqV'�'����(K>ɨCN*��
���G`>^�X�`���K:��K,��xA	�`���#0�=Y��X�`��+w�ÏT�X�X�`���+���k,��x���8X�`���+����,����1���ogЯg���IՏ�V?X>��R>�����G`>^��X�`����'���,��x�'�`���#0/Y�,_�|�㕪`������|�P�}
X�`���K{���,����:o����˷\�.\�j��ţ?OC���@,_<X�x�|����W����/X>���w�����G`>^��X�`��Ǖ���,���I�����˷,�!��H_��	`���#0�� ��~�|��`������|\G�?�|����ˈ���^b�^c�/,_X�`��gO��@��/X�e�a!��\�v?X�`���Un���,���>�`���#0����/�����|\��?�|��������/X>�ٓ�V����oY�KX���ӟV?�~�|��Y`�������O��V?X>�q�2�����G`>.��X�`��������,�����X�`�������,���� �`���+|����Inl>/������l�檈�bƳ�" �8�yU�$����nl>������D��`��»a�I�����a�1������[��o�}�����[lٸ� ���<In}G�??{��}���E���{韷�?/��[n��S�Wv����S��J��eW/��Ot�^8�-��{mߎuY��&�H&P_���k���'��P��4��𯯏�Y�ׇܮh|C�<�j�8�����Xumo�#�מ�|�ڳ��_{V�KӍ��];�����DSu���bo5�E����d+����VF��k�q�al�t��6uR��`J��}�ض�p�Y�ׯ=����g5_��чƹ����ܦة��L�&W�c�p�ڳ��_{V��k�ʷdc�2llS�UJ���hmtD�� ��|>���d�6q�e�4F�����1��4~Dmy1�f4��i3��Ç����}֗�r�e9z3�>ֶ)]�������Y���n���0�)]T)q�ƚ6�e)�}�t�g5_�/ʒ�X3�<B4mA��i�\�Xji��׳�_eڒ�*K3�0�!2���J��4}���l�K������uj�&C����f'Eӛt�[�.��~,�pi��j>��_����}����q���d-���N�۽���MY	C24%:Ȑ�AC2d��%�d�eH2T�V��(��
��@��<�d(�
!Q�"�P>��C24�{Ph.k��6,o�C�7�27�R7ʒ����`ٛ`�`��`	ei�u��qX'XGY���,�;Xw�<�`yei*�	�q����Q��������}	f�N��@L�<�@ٗ`���"
���nʾTW]+͙ KS�,P~:X�E�V��	��Q����	�$�(��=,��,q,,���P���1�\0YrM�*/d��q�%.*c����a8�W��1��x��q�%����(KS-P.8XrUS׍�	��Q����	6��8��r�1��x��q�%.9��(K��bP.8X�����L�<�����aL��x���Q�x]3�	��#,��,��[,�GXGY�u�0&X/`�q�%^�c���X_��}��|�+���au�t.Y��+��Ϭ�����_1~�/���U��TX�~�,n�WVRa��y��U�_5XI�5�.�΋�`<��J*�i���y��4XI�5�QT�:/���+������*Я�t�U>Ϛ�	��u^,�VRa��y� �U�_5XI���	�:�K��th��f�*�.%٥��HGx���R���g:�tԗ
-���7�:��Q`*��C�����VG��В-�a��S�%Z^���[5�BK�ic�� #E�BK:��6FǷ:�L��thy��΋]�BK:��VIǷ:�L��thy͕�o�ވ)���eNG�9]�BK:��NǷ:�L��thy-��out�
-���D���2Zҡ嵕:���e*��C�kDu|���ThI��׺��VG��В-����0IG��В-�=��.S�%Z^C��[]�BK�i��+}�������:����2���ThI������VG��В-���.S�%Z����[]�BK:�\�AǷ:�L��th�v��out�
-�������.:�L��th����out�
-��rM���2Zҡ��.:���e*��C�5jt|���Li)��.:�,��2Zҡ�A:���e*�t�0��eAG��В-�p��.S�%Z�E��[]�BK:�\SKŷQG��В-���.S�%Z�q��[]�BK:�\�MǷ:�L������`QG�E]�BK:�\;OǷJU>��|�貨�ˢ�.S�%Z�e��[]�BK:�\�QǷ:�L��th����out�
-��r�L�:�L��th�֧�out�
-��r�R���2Zʣ}�#����6��ʛ*��u7T�PT}���a�he�6�F++�d7ZY����Ty{Y�u��x^�m��R�z���z���T��he���֨/&z�6}�j�k[�n5�R�}�L��9��&��v�ܚ��F,6h�jf���/[�LQ��Fj��)��;�m5��⵽ ����x��V3%�L�1SC�xL.^�=��L;�e��49�d���˾6i���U�}V�e�ruXȲruT���1�ɩ�6!��i��;�U��6����,+W��e�_��d��M[�v4u�	����3>v��:j��Yp���yD���iD���~�q�al�t'�uuR��`J��}�ض��,+W��e�_��\���C�\h�sm�bS��CM�o��ӏ1R��,+W��e�_��-�X%M�d%EN�R�qu5ZQg�_Q���W�e%#c�Ml��6I�PPcZ�4��C�dt�і9c@���1 ���+
�O�.�;�/+~���7��cm�ҥ\��,+W�(���+��q,�:c�Ч,U�|�k�P�U���1#�dY�zEEYR�`�`S�M[�hz�4c���x�%�����-���4#C�c�.�J��4}���l���2YV���Pۑ���}LS���MJ,֤+-��K;d��YV�Y~����O���{�˫���1������y̷}7#��C��2*�d�N�0�d�NO� D Cvzz!�ӓHȐ��jB�@���B2d���"�!{xr�I����K۰�M�č�d�1L��M�䍲d��1L��M���d�1L�N�$��d�0L�<�`ye�^�`�p�o���,��,���,�;XGY��7Q&Xw�<��d��0L�<�`ye���a�8,�{XGY�w0&ܓܣX��<�����`L�<�aye��a��`y���8��_�1��x��q�%��c��� ��(K\_Ƅ{&�{(����Q���	��,��,q�	,�XGY�:�W?�<aye���Ø`y<��8���1��n�^o��x��q�%^oc�����(K�����,��,�zB,��<�fi�����S���>�URa%V�_�;E[�U��TX�~��m�WVRa��E �U�_5XI�5�.�.J A<��J*�i���E��4XI�5�QT��(��+�������*Я���j���?h�@�j��
��/�������J*��M��0�Q\*��C��6��VIu)�.�E:t��
-����:��Q_*��C�����VG��В-���[�BK:���AǷ:JL��thy-��ouԘ
-�����(2Zҡ�1:��Qe*��C�k|t^,��2Zҡ�J:���e*��C�k�t|��FL镘�.s:����2Zҡ�5p:���e*��C�k�t|���ThI���$��VG��В-����.S�%Z^#��[]�BK:���UǷ:�L��thyͮ·I:�L��thy�out�
-���j���2Zҡ��:�U�ZQ�sE]�ut���e*��C�k�u|���ThI��k��VG��В-�J��.S�%Z����[]�BK:�\�BǷ:�L��th���o��.S�%Z�%��[]�BK:�\EǷ:�L��th����out�
-��r��*�$SZJ��˂�.:�L��th�f��out�
-��r�#���2Zҡ�N:���e*��C˵�t|���ThI��kj��6��2Zҡ��`:���e*��C�5�t|���ThI��k���VG��В-ל��.S�%Z����[�*Je>ttY��eQG��В-�2��.S�%Z�ɨ�[]�BK:�\[RǷ:�L��th�F��o]�BK:�\�SǷ:�L��th�f��out�
-�Ѿn]����X�ڏ�	m�Mg���f(��vk�0o��R�v���j������he���F++��7ZY�n���J=�VV*Ho��R�ykԁ��k��n5��ߵ�U���D���[�`bxm�Эf0Q���V3����]*���D��^�[�`�xm�ŭf0Q�����Q�k���iǺ��h��(�	��.�ڤISOTW�.��YM���*�����+��P'��ڄ0���Bo�8V]������_��\�K���~ɲ��g��v�h�:bM�yg|�:��u�9��+8�JFΰr�/64�m��D���nC�:LI��/۶���e�_��\�K���~}h��q�MVl
�z���m�v�1F
���e�_��\�U�%��)c���ȩR�1��Fk�#���+ʲr����dd̶��-S�&�
jL��T~蓌�4�2gȰ�1dX�zEa�)��t'�e�O ��r�fp}�mS���W�e��eY�zEU7�Ygl������|cMʲ��>f�,+W��(Kjb�l��iMOc��RK�u�,+��ƶ$��Ҍ4i��}��*][��]���2��dY���CmG�*S�1MɊ�7)�X����~,�16fY9f��M�Ͽ��xx�����{G������i��}����~�����w�~+yf6{�,y ���ooneO�f�OH�o U�`J(9ͼ�G�y=K!�zg^�L�7P�Ҿ�2�,��/š ��B����?�}�8y��BF��>^F��Ko@+#H�`ei^�C�#���u��	2��i��kE�p�?'������|]��OCu�sy��)s}�2E~z�K��7������	��f��=Ü}٩������{R0&���P���
.k TRu��0���PH�&L���K'����������! �A�v��A�xZ�c���1���� *�P��>�B��1bٟ0v�~���?=7�������`~����x����"	j~׸��H���WB
���WB
�	;}/#������B
�	;}�oO�'��D9T!w�؄��\�dP����Fl�Nk�b��Vb�C�0�!R-"���xc��h @�%@��۰��$R@�3)�br0��܆=����'� y� �Xn��H9 �؝���g6�\� �Xn�� ���X�\� �Xn��DI9 �؉'l�ê,) �:q�$�{X&� d�ia��]L�ǟp���nmfR8d�1�HH	H�r����T�X��= �m��; @.���n�>�MN�&��3&�43���3� ̚����_� �� ��r�����$|�79��[�>�=gR$�V?�Oy< ��r\��S@.����� @.�gf��ǥp��+�I�3�s&E �6��O�6��2�0���9����p rq�b���
� ����r\O���`^,��u*�yqȧK�kK.j����?��-V�,��\�ά�>_��E�R�weK�������Jq� �������C��A���#0_R2`�-�~^/���|i���b{��b�̗f	`�-�p^/���|v�حg�?,�b����_�b��;;3/�G`>�_l�����|�y(z>��+`BB�h�E	\��e	�u�|U�����dI8Z��h�Bh�&$4!���!Z��		M��n�}��,`BB��h�u��Є���	Ƈh�&\q��H�������Є�8�C����V��j�U��Є�
�C���О�����z�~嚊����7h��U��Є�r�C����W=�}�V1`BB�-��*LHhB^m��!Zŀ		M�+��>D�0!�	y�ڇh�&$4!�ADL��-`BB�
I�ѲLHhB{R��C�l.�^^|��߉�?�)��--[<Z��		M���>D�0!�	yq3ڇh�&$4!/�F�-[���&��h�e��Є��R0Ƈh�&\G�\a�Z�����k�}�V1`BBr]��*LHhB���!Z��		M�'�>��q�/rA˖��--[���&�'�`|��-`���+�����	h&$4!�TA��b���&�r0h�U��Є\��È�-`BBr��ѲLHhB.��!Z��		MhO�4��-[���m�.���h�*LHhB�$��!|�>|�>Z�D���h&$4!W�B�-[���&��ch�e��Є\9�C�l�����}X�e��Є\��C�l����}��-`B�F�q��E�ō��n�)l�����������Xzf�0ɖ�����/�nl��S����������4>���m5 ����u[,� o5 ��.n[Hq�o��͡/W�޾������7l������/�"�՞4��{um5���Ŋ<~f�CQDTK{�-���U���u�����P�ڱ.�2�4ىd���˾6i��U�i���^��/Y�/�]��>�:���&�q4mzcǱ���&o֗�?�����j����_	��v�h�:bM�yg|�:�}�=�py�����\ ��ũ@F��o�@��V��q)~�6�����]���m{����_�����?����}h��q�M�m
�z���m�g�1F
��?�����j����-�X%���>EB�R�qu5ZQg/�g������b�j�8�2uX����ƴ�iL�>I�H�-/�ߌ��oF��a�)�t��e��95-Go���6�K��ğ��V��U7�Ygl��?��I|cMʲ��>^����_�/ʒ�X3��B4mA��i�\�Xji�����_ڒ�*K3�0��3�	�JW�4}���l���*��_��>�v��2u��hz�n|k�u]׏�.�?Y���7��vw���a�>����˙F��}��=Oƹ�/�g�U���<O�x���P��N��N�N��MMK
����Ц�����Ǥ�����[8nḅ��[8nḅ�ij���]�$h�����6�v�6���6�(N~������rR�QNZ4�I��R�����A��y� �~:j��[�~x�;i�r7ϟ�&�G��W
���K8:����Q�Ly�jc	�N��#�dQ�|��|$*�����$RB��E��QH�>���ZB�(�e�`�*��*zDW�!��D"�g�jiX�|T,��J�D۬��P"By�v�����i?w���4�G����V�K(iz�����D������|�P�ރ�Z�r�ΒP��h۹��KBY�����dK"Y��Y�nͶ r��O�;a���%�,��,{l�w$����>��7��u���o�n������͎ЧC�<�>r�C��!�<>
�C�ӡ�<T|:T,����CէC��P��P�8D/ޠ�;�;�����!��Zz�^<BK�ЋKh�z�	-�B/N��W��+�t����~q/~qK�����H1׼�?�����a����o����r��|�8��t�>�_؛@'���b�~���+_�~�3��G��b~�~���Ç���n������ŷrr������ɑ��O�3}��K��#���٩�����t��_O?>���Lvw����Ӑ>��{�k���8��ǻǡ߽{NW�:�����t���K ǧ�<��� $	�������C�÷ɝ�m���&��19���%5�9߷1XoR�XS�3�ƺ�T�O�)c�iw�O��}wh��������.�Vs`�}��~��=v�O���|�yCU"b���{t�WGG|y|$	�G��W�P���#���?>�A�"�`��駒��'���1wr��������N�'��ɱ�2?�D���U��:9V��'���1����S�߻�o�?�w�}Ko�[�r����?�)B��O)����7���ۿ�Ꮯ3�e�����Y>ݢ�{�����~��8P�GS�C��ʻICi��2eض������n!�~u�##�����TLq2�tt��_N�=���D�\���a@OY��r≦�����C�p:)��yE�vh������V���p���R2'����"b�L,��:���ߣ�7�2��t�k@� �GY��(��s���яܙ��>�y�������*�z�O��?߿���i��F����/��~�r$ڣ���Qg��b�OCQ/��H�Z�����~Sw]�$��}���X�zl}�L��C�ʑ�]�����>�g�y�9J\��:l����Ί�w�_T�OK3�P�¾L�茵Ȏv�:���t�q�ѵ�������h7��E��X0]��ӳ.�u�#���?EĹ����j��IW����X'��}8wKW���8t���K>N�i���ٿ��W����o�wUY��;�`Y9]�JO���|ր�D���߾6�,�����>]|�F�~KE]�7��޺ڽ>{<�����ԓ��8��|����8ڡ��+��V�$����˙�M��|X���A�����i��	d���J�T�8���2#N���" x(��6�;�{t ���C�|'.���FI�7�Q�ӊp���&a�YΜ�{� B'��ڡ��uuF����z�L3a��ۇ���2�ɽ;C.�N$��k�]^��]��#�p/�1�/�~��O-����7�۩}^��t?�?~k�������?�?��ԓӼ���Rx�x�n���?}�7�n��Q����w���O�n�h|26��gLI�e�L?6?�DM���퇇��篛�'ۿ|��w;~����|���.~�߾���yx���Q֞�x�l��xs�4oWN�+�}��w�_S(�F���Q�Q���~�Q1*^h7G?Iψ��Ӓ�ˉ��i7G�K.��Qn
�WZ���5������q}k�L/�_�5��Q2;�v?9h���� )��ෆ��j�z�N��!�M�[� RH�ෆ@�J�F��0 6��*8�p~c PN��M�_�V��/M7�~���x��oc�<���1~vZ8?����|����W���/d�X)�7��mS�"o��uvZ�~>��ho92����On�M�Ue�L5��r%�T��d�8d2*�>�dTܖ��rѬ�W��L���r^f�P]u-<b�s˪oŠ��ͭ��{oo�-����E_��}�p��%|�����M~��Z�����<��?�S����:<پ��}�#��Y_���I�-� U��y���l���!K"����p�'`�R���l(�������:�g 7��E�z��Y��0QxR~~�L ����/&�	Ƭތ��!������Cփ,_�p��H�0��Q�r>L��o�uĜ<���
�o&t9L6W^�
�i�a{9,n���bZy�������Y�+���ǿ�?��z[�s��Ϸr��|檦�p�^�6��ҋ�4ʁ�����EN4��2.�|wV��8�<o5��x�-���iS�ʃ���$~s�6�8M�vp�:�$�|��ͳ���+y������V��̧��2��u[u�8E��R{�Ȝ�8��g�#��f���s+y2��i�y��3�����8����PK   WlKTzײ�+*  ��            ��    cirkitFile.jsonPK      =   X*    